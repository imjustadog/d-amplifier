library verilog;
use verilog.vl_types.all;
entity verilog_yunfang_vlg_tst is
end verilog_yunfang_vlg_tst;
